// F12 verilog III
// Course   : HE1026 Digital teknik
// Datum    : 2025-11-25

module top(input [8:1] GP, input GP9, input GP18, output [8:1] LED)
    //

endmodule
